* Top cell name: cnt_control

.SUBCKT nand2 in0 in1 out vdd vss
    Mm1 net9 in1 vss vss n_mos l=30n w=200n m=1 nf=1
    Mm0 out in0 net9 vss n_mos l=30n w=200n m=1 nf=1
    Mm3 out in1 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm2 out in0 vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT nand3_r in0 in1 in2 out rst vdd vss
    Mm3 out rst vss vss n_mos l=30n w=300n m=1 nf=1
    Mm2 net6 in2 vss vss n_mos l=30n w=300n m=1 nf=1
    Mm1 net7 in1 net6 vss n_mos l=30n w=300n m=1 nf=1
    Mm0 out in0 net7 vss n_mos l=30n w=300n m=1 nf=1
    Mm7 net21 rst vdd vdd p_mos l=30n w=200n m=1 nf=1
    Mm6 out in2 net21 vdd p_mos l=30n w=200n m=1 nf=1
    Mm5 out in1 net21 vdd p_mos l=30n w=200n m=1 nf=1
    Mm4 out in0 net21 vdd p_mos l=30n w=200n m=1 nf=1
.ENDS

.SUBCKT nand3 in0 in1 in2 out vdd vss
    Mm4 net016 in2 vss vss n_mos l=30n w=300n m=1 nf=1
    Mm1 net3 in1 net016 vss n_mos l=30n w=300n m=1 nf=1
    Mm0 out in0 net3 vss n_mos l=30n w=300n m=1 nf=1
    Mm5 out in2 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm3 out in1 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm2 out in0 vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT dff_st_ar clk d q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi3 n1 d n3 vdd vss nand2
    Xi2 n3 n0 n2 vdd vss nand2
    Xi6 clk n0 n3 n1 rst vdd vss nand3_r
    Xi7 clk n2 rst' n0 vdd vss nand3
.ENDS

.SUBCKT nor5 in0 in1 in2 in3 in4 out vdd vss
    Mm4 out in4 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm3 out in0 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm2 out in1 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm1 out in3 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm0 out in2 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm9 net12 in4 vdd vdd p_mos l=30n w=400n m=1 nf=1
    Mm8 net13 in3 net12 vdd p_mos l=30n w=400n m=1 nf=1
    Mm7 net14 in2 net13 vdd p_mos l=30n w=400n m=1 nf=1
    Mm6 net15 in1 net14 vdd p_mos l=30n w=400n m=1 nf=1
    Mm5 out in0 net15 vdd p_mos l=30n w=400n m=1 nf=1
.ENDS

.SUBCKT inv in out vdd vss
    Mm0 out in vss vss n_mos l=30n w=100n m=1 nf=1
    Mm1 out in vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT nor2 in0 in1 out vdd vss
    Mm1 out in1 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm0 out in0 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm3 net5 in1 vdd vdd p_mos l=30n w=200n m=1 nf=1
    Mm2 out in0 net5 vdd p_mos l=30n w=200n m=1 nf=1
.ENDS

.SUBCKT nor4 in0 in1 in2 in3 out vdd vss
    Mm3 out in3 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm2 out in2 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm1 out in1 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm0 out in0 vss vss n_mos l=30n w=100n m=1 nf=1
    Mm7 net24 in3 vdd vdd p_mos l=30n w=400n m=1 nf=1
    Mm6 net23 in2 net24 vdd p_mos l=30n w=400n m=1 nf=1
    Mm5 net25 in1 net23 vdd p_mos l=30n w=400n m=1 nf=1
    Mm4 out in0 net25 vdd p_mos l=30n w=400n m=1 nf=1
.ENDS

.SUBCKT nand5 in0 in1 in2 in3 in4 out vdd vss
    Mm4 net21 in4 vss vss n_mos l=30n w=400n m=1 nf=1
    Mm3 net22 in3 net21 vss n_mos l=30n w=400n m=1 nf=1
    Mm2 net23 in2 net22 vss n_mos l=30n w=400n m=1 nf=1
    Mm1 net24 in1 net23 vss n_mos l=30n w=400n m=1 nf=1
    Mm0 out in0 net24 vss n_mos l=30n w=400n m=1 nf=1
    Mm9 out in0 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm8 out in4 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm7 out in3 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm6 out in1 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm5 out in2 vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT cnt_rst_fb cnt_data<0> cnt_data<1> cnt_data<2> cnt_data<3> cnt_data<4> cnt_data<5>
                   + cnt_data<6> cnt_data<7> cnt_data<8> cnt_data<9> cnt_data<10> cnt_data<11>
                   + cnt_data<12> cnt_data<13> cnt_data<14> extclk_cnt<0> extclk_cnt<1>
                   + extclk_cnt<2> extclk_cnt<3> extclk_cnt<4> out out' ready2 vdd vdl_rst vss
    Xi7 cnt_data<12> cnt_data<13> cnt_data<14> vdl_rst ready2 net44 vdd vss nor5
    Xi0 extclk_cnt<0> extclk_cnt<1> extclk_cnt<2> extclk_cnt<3> extclk_cnt<4> net48 vdd vss nor5
    Xi4 cnt_data<8> cnt_data<9> cnt_data<10> cnt_data<11> net45 vdd vss nor4
    Xi3 cnt_data<4> cnt_data<5> cnt_data<6> cnt_data<7> net27 vdd vss nor4
    Xi2 cnt_data<0> cnt_data<1> cnt_data<2> cnt_data<3> net34 vdd vss nor4
    Xi5 net48 net34 net27 net45 net44 out' vdd vss nand5
    Xi8 out' out vdd vss inv
.ENDS

.SUBCKT nand4 in0 in1 in2 in3 out vdd vss
    Mm3 net17 in3 vss vss n_mos l=30n w=400n m=1 nf=1
    Mm2 net18 in2 net17 vss n_mos l=30n w=400n m=1 nf=1
    Mm1 net19 in1 net18 vss n_mos l=30n w=400n m=1 nf=1
    Mm0 out in0 net19 vss n_mos l=30n w=400n m=1 nf=1
    Mm7 out in0 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm6 out in3 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm5 out in2 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm4 out in1 vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT cnt_vdl_rst_fb cnt_data<0> cnt_data<1> cnt_data<2> cnt_data<3> cnt_data<4> cnt_data<5>
                       + cnt_data<6> cnt_data<7> cnt_data<8> cnt_data<9> cnt_data<10> cnt_data<11>
                       + cnt_data<12> cnt_data<13> cnt_data<14> out ready_clk vdd vss
    Xi3 cnt_data<12> cnt_data<13> cnt_data<14> ready_clk net1 vdd vss nor4
    Xi2 cnt_data<8> cnt_data<9> cnt_data<10> cnt_data<11> net8 vdd vss nor4
    Xi1 cnt_data<4> cnt_data<5> cnt_data<6> cnt_data<7> net034 vdd vss nor4
    Xi0 cnt_data<0> cnt_data<1> cnt_data<2> cnt_data<3> net035 vdd vss nor4
    Xi4 net035 net034 net8 net1 net031 vdd vss nand4
    Xi5 net031 out vdd vss inv
.ENDS

.SUBCKT inv_dh in out vdd vss
    Mm0 out in vss vss n_mos l=30n w=200n m=1 nf=1
    Mm1 out in vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT dff_st_ar_dh clk q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi2 n3 n0 n2 vdd vss nand2
    Xi6 clk n0 n3 n1 rst vdd vss nand3_r
    Xi7 clk n2 rst' n0 vdd vss nand3
    Xi8 n1 n3 vdd vss inv_dh
.ENDS

.SUBCKT cnt_control cnt_data<0> cnt_data<1> cnt_data<2> cnt_data<3> cnt_data<4> cnt_data<5>
                    + cnt_data<6> cnt_data<7> cnt_data<8> cnt_data<9> cnt_data<10> cnt_data<11>
                    + cnt_data<12> cnt_data<13> cnt_data<14> cnt_ready cnt_rst cnt_rst'
                    + extclk_cnt<0> extclk_cnt<1> extclk_cnt<2> extclk_cnt<3> extclk_cnt<4> ext_clk
                    + ready_clk rst_glob rst_glob' vdd vdl_rst_loc vdl_rst_loc' vss
    Xi10 pre_rst vdl_rst_loc vdl_rst_rst_loc vdl_rst_rst_loc' vdl_rst_loc' vdl_rst_loc vdd vss
         + dff_st_ar
    Xi8 ready_clk net019 vdl_rst_0 vdl_rst_0' vdl_rst_rst vdl_rst_rst' vdd vss dff_st_ar
    Xi1 ready_clk ready2 cnt_ready vdl_rst_1' cnt_rst_pre cnt_rst_pre' vdd vss dff_st_ar
    Xi0 ext_clk net19 cnt_rst_loc cnt_rst_loc' cnt_rst_rst cnt_rst_rst' vdd vss dff_st_ar
    Xi2 extclk_cnt<0> extclk_cnt<1> extclk_cnt<2> extclk_cnt<3> net27 net19 vdd vss nor5
    Xi9 ready2 net019 vdd vss inv
    Xi3 extclk_cnt<4> net27 vdd vss inv
    Xi14 vdl_rst_0' vdl_rst_1' vdl_rst_loc vdd vss nand2
    Xi17 vdl_rst_0' cnt_rst_pre' cnt_rst vdd vss nand2
    Xi11 cnt_rst_pre' vdl_rst_rst_loc' vdl_rst_rst vdd vss nand2
    Xi5 cnt_rst_loc' rst_glob' cnt_rst_pre vdd vss nand2
    Xi18 vdl_rst_0 cnt_rst_pre cnt_rst' vdd vss nor2
    Xi15 vdl_rst_0 cnt_ready vdl_rst_loc' vdd vss nor2
    Xi12 cnt_rst_pre vdl_rst_rst_loc vdl_rst_rst' vdd vss nor2
    Xi6 cnt_rst_loc rst_glob cnt_rst_pre' vdd vss nor2
    Xi7 cnt_data<0> cnt_data<1> cnt_data<2> cnt_data<3> cnt_data<4> cnt_data<5> cnt_data<6>
        + cnt_data<7> cnt_data<8> cnt_data<9> cnt_data<10> cnt_data<11> cnt_data<12> cnt_data<13>
        + cnt_data<14> extclk_cnt<0> extclk_cnt<1> extclk_cnt<2> extclk_cnt<3> extclk_cnt<4>
        + cnt_rst_rst cnt_rst_rst' ready2 vdd vdl_rst_loc vss cnt_rst_fb
    Xi16 cnt_data<0> cnt_data<1> cnt_data<2> cnt_data<3> cnt_data<4> cnt_data<5> cnt_data<6>
         + cnt_data<7> cnt_data<8> cnt_data<9> cnt_data<10> cnt_data<11> cnt_data<12> cnt_data<13>
         + cnt_data<14> pre_rst ready_clk vdd vss cnt_vdl_rst_fb
    Xi4 ready_clk ready2 net03 cnt_rst_pre cnt_rst_pre' vdd vss dff_st_ar_dh
.ENDS
