* Top cell name: core_control

.SUBCKT nand2 in0 in1 out vdd vss
    Mm1 net9 in1 vss vss n_mos l=30n w=200n m=1 nf=1
    Mm0 out in0 net9 vss n_mos l=30n w=200n m=1 nf=1
    Mm3 out in1 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm2 out in0 vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT inv in out vdd vss
    Mm0 out in vss vss n_mos l=30n w=100n m=1 nf=1
    Mm1 out in vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT mux2 in0 in1 out sel vdd vss
    Xi2 in0 net7 net9 vdd vss nand2
    Xi1 in1 sel net10 vdd vss nand2
    Xi0 net10 net9 out vdd vss nand2
    Xi3 sel net7 vdd vss inv
.ENDS

.SUBCKT mux4 in<0> in<1> in<2> in<3> out sel<0> sel<1> vdd vss
    Xi2 in<2> in<3> net5 sel<0> vdd vss mux2
    Xi1 in<0> in<1> net6 sel<0> vdd vss mux2
    Xi0 net6 net5 out sel<1> vdd vss mux2
.ENDS

.SUBCKT nand3_r in0 in1 in2 out rst vdd vss
    Mm3 out rst vss vss n_mos l=30n w=300n m=1 nf=1
    Mm2 net6 in2 vss vss n_mos l=30n w=300n m=1 nf=1
    Mm1 net7 in1 net6 vss n_mos l=30n w=300n m=1 nf=1
    Mm0 out in0 net7 vss n_mos l=30n w=300n m=1 nf=1
    Mm7 net21 rst vdd vdd p_mos l=30n w=200n m=1 nf=1
    Mm6 out in2 net21 vdd p_mos l=30n w=200n m=1 nf=1
    Mm5 out in1 net21 vdd p_mos l=30n w=200n m=1 nf=1
    Mm4 out in0 net21 vdd p_mos l=30n w=200n m=1 nf=1
.ENDS

.SUBCKT nand3 in0 in1 in2 out vdd vss
    Mm4 net016 in2 vss vss n_mos l=30n w=300n m=1 nf=1
    Mm1 net3 in1 net016 vss n_mos l=30n w=300n m=1 nf=1
    Mm0 out in0 net3 vss n_mos l=30n w=300n m=1 nf=1
    Mm5 out in2 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm3 out in1 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm2 out in0 vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT dff_st_ar clk d q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi3 n1 d n3 vdd vss nand2
    Xi2 n3 n0 n2 vdd vss nand2
    Xi6 clk n0 n3 n1 rst vdd vss nand3_r
    Xi7 clk n2 rst' n0 vdd vss nand3
.ENDS

.SUBCKT tff_st_ar clk q q' rst rst' vdd vss
    Xi8 clk q' q q' rst rst' vdd vss dff_st_ar
.ENDS

.SUBCKT freq_scaler in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> rst rst' vdd vss
    Xi11 out<6> out<7> net32 rst rst' vdd vss tff_st_ar
    Xi10 out<5> out<6> net34 rst rst' vdd vss tff_st_ar
    Xi9 out<4> out<5> net35 rst rst' vdd vss tff_st_ar
    Xi8 out<3> out<4> net36 rst rst' vdd vss tff_st_ar
    Xi7 out<2> out<3> net37 rst rst' vdd vss tff_st_ar
    Xi6 out<1> out<2> net38 rst rst' vdd vss tff_st_ar
    Xi5 out<0> out<1> net39 rst rst' vdd vss tff_st_ar
    Xi4 net16 out<0> net40 rst rst' vdd vss tff_st_ar
    Xi3 net14 net16 net41 rst rst' vdd vss tff_st_ar
    Xi2 net12 net14 net42 rst rst' vdd vss tff_st_ar
    Xi1 in net12 net43 rst rst' vdd vss tff_st_ar
.ENDS

.SUBCKT mux8 in<0> in<1> in<2> in<3> in<4> in<5> in<6> in<7> out sel<0> sel<1> sel<2> vdd vss
    Xi1 in<4> in<5> in<6> in<7> net4 sel<0> sel<1> vdd vss mux4
    Xi0 in<0> in<1> in<2> in<3> net5 sel<0> sel<1> vdd vss mux4
    Xi2 net5 net4 out sel<2> vdd vss mux2
.ENDS

.SUBCKT core_control conf_rochoose<0> conf_rochoose<1> conf_roen conf_rofreq<0> conf_rofreq<1>
                     + conf_rofreq<2> conf_rst conf_rst' ext_rst ext_rst' ro_in<0> ro_in<1> ro_in<2>
                     + ro_in<3> ro_out vdd vss
    Xi0 ro_in<0> ro_in<1> ro_in<2> ro_in<3> net1 conf_rochoose<0> conf_rochoose<1> vdd vss mux4
    Xi1 net07 net08<0> net08<1> net08<2> net08<3> net08<4> net08<5> net08<6> net08<7> ext_rst
        + ext_rst' vdd vss freq_scaler
    Xi2 net08<0> net08<1> net08<2> net08<3> net08<4> net08<5> net08<6> net08<7> ro_out
        + conf_rofreq<0> conf_rofreq<1> conf_rofreq<2> vdd vss mux8
    Xi3 net1 conf_roen net07 vdd vss nand2
    Xi5 ext_rst ext_rst' vdd vss inv
    Xi4 conf_rst conf_rst' vdd vss inv
.ENDS
