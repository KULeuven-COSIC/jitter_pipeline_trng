* Top cell name: vdl_oo_3

.SUBCKT inv_oo_dc_0 in out vdd vss
    Mm0 out in vss vss n_mos l=30n w=100n m=1 nf=1
    Mm1 out in vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT inv_oo_dc_1 conf conf' in out vdd vss
    Mm1 net7 conf vss vss n_mos l=30n w=100n m=1 nf=1
    Mm0 out in net7 vss n_mos l=30n w=100n m=1 nf=1
    Mm3 net5 conf' vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm2 out in net5 vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT vdl_oo_2 conf'<0> conf'<1> conf'<2> conf'<3> conf'<4> conf'<5> conf'<6> conf'<7> conf'<8>
                 + conf'<9> conf'<10> conf'<11> conf'<12> conf'<13> conf'<14> conf'<15> conf<0>
                 + conf<1> conf<2> conf<3> conf<4> conf<5> conf<6> conf<7> conf<8> conf<9> conf<10>
                 + conf<11> conf<12> conf<13> conf<14> conf<15> in out vdd vss
    Xi1 int out vdd vss inv_oo_dc_0
    Xi0 in int vdd vss inv_oo_dc_0
    Xi17 conf<15> conf'<15> int out vdd vss inv_oo_dc_1
    Xi16 conf<7> conf'<7> in int vdd vss inv_oo_dc_1
    Xi15 conf<14> conf'<14> int out vdd vss inv_oo_dc_1
    Xi14 conf<6> conf'<6> in int vdd vss inv_oo_dc_1
    Xi13 conf<13> conf'<13> int out vdd vss inv_oo_dc_1
    Xi12 conf<5> conf'<5> in int vdd vss inv_oo_dc_1
    Xi11 conf<12> conf'<12> int out vdd vss inv_oo_dc_1
    Xi10 conf<4> conf'<4> in int vdd vss inv_oo_dc_1
    Xi9 conf<11> conf'<11> int out vdd vss inv_oo_dc_1
    Xi8 conf<3> conf'<3> in int vdd vss inv_oo_dc_1
    Xi7 conf<10> conf'<10> int out vdd vss inv_oo_dc_1
    Xi6 conf<2> conf'<2> in int vdd vss inv_oo_dc_1
    Xi5 conf<9> conf'<9> int out vdd vss inv_oo_dc_1
    Xi4 conf<1> conf'<1> in int vdd vss inv_oo_dc_1
    Xi3 conf<8> conf'<8> int out vdd vss inv_oo_dc_1
    Xi2 conf<0> conf'<0> in int vdd vss inv_oo_dc_1
.ENDS

.SUBCKT nand2_dnw in0 in1 out vdd vss
    Mm0 out in0 net9 vss n_mos l=30n w=200n m=1 nf=1
    Mm1 net9 in1 vss vss n_mos l=30n w=200n m=1 nf=1
    Mm3 out in1 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm2 out in0 vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT vdl_oo_3 conf'<0> conf'<1> conf'<2> conf'<3> conf'<4> conf'<5> conf'<6> conf'<7> conf'<8>
                 + conf'<9> conf'<10> conf'<11> conf'<12> conf'<13> conf'<14> conf'<15> conf<0>
                 + conf<1> conf<2> conf<3> conf<4> conf<5> conf<6> conf<7> conf<8> conf<9> conf<10>
                 + conf<11> conf<12> conf<13> conf<14> conf<15> enable out vdd vss
    Xi0 conf'<0> conf'<1> conf'<2> conf'<3> conf'<4> conf'<5> conf'<6> conf'<7> conf'<8> conf'<9>
        + conf'<10> conf'<11> conf'<12> conf'<13> conf'<14> conf'<15> conf<0> conf<1> conf<2>
        + conf<3> conf<4> conf<5> conf<6> conf<7> conf<8> conf<9> conf<10> conf<11> conf<12>
        + conf<13> conf<14> conf<15> nand out vdd vss vdl_oo_2
    Xi1 out enable nand vdd vss nand2_dnw
.ENDS
