* Top cell name: cnt_data_chain

.SUBCKT nand2 in0 in1 out vdd vss
    Mm1 net9 in1 vss vss n_mos l=30n w=200n m=1 nf=1
    Mm0 out in0 net9 vss n_mos l=30n w=200n m=1 nf=1
    Mm3 out in1 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm2 out in0 vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT nand3_r in0 in1 in2 out rst vdd vss
    Mm3 out rst vss vss n_mos l=30n w=300n m=1 nf=1
    Mm2 net6 in2 vss vss n_mos l=30n w=300n m=1 nf=1
    Mm1 net7 in1 net6 vss n_mos l=30n w=300n m=1 nf=1
    Mm0 out in0 net7 vss n_mos l=30n w=300n m=1 nf=1
    Mm7 net21 rst vdd vdd p_mos l=30n w=200n m=1 nf=1
    Mm6 out in2 net21 vdd p_mos l=30n w=200n m=1 nf=1
    Mm5 out in1 net21 vdd p_mos l=30n w=200n m=1 nf=1
    Mm4 out in0 net21 vdd p_mos l=30n w=200n m=1 nf=1
.ENDS

.SUBCKT nand3 in0 in1 in2 out vdd vss
    Mm4 net016 in2 vss vss n_mos l=30n w=300n m=1 nf=1
    Mm1 net3 in1 net016 vss n_mos l=30n w=300n m=1 nf=1
    Mm0 out in0 net3 vss n_mos l=30n w=300n m=1 nf=1
    Mm5 out in2 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm3 out in1 vdd vdd p_mos l=30n w=100n m=1 nf=1
    Mm2 out in0 vdd vdd p_mos l=30n w=100n m=1 nf=1
.ENDS

.SUBCKT dff_st_ar clk d q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi3 n1 d n3 vdd vss nand2
    Xi2 n3 n0 n2 vdd vss nand2
    Xi6 clk n0 n3 n1 rst vdd vss nand3_r
    Xi7 clk n2 rst' n0 vdd vss nand3
.ENDS

.SUBCKT tff_st_ar clk q q' rst rst' vdd vss
    Xi8 clk q' q q' rst rst' vdd vss dff_st_ar
.ENDS

.SUBCKT cnt_data_chain out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> out<8> out<9> out<10> out<11> out<12> out<13> out<14> rand_in rst rst' vdd vss
    Xi15 out<13> out<14> net10 rst rst' vdd vss tff_st_ar
    Xi14 out<12> out<13> net17 rst rst' vdd vss tff_st_ar
    Xi13 out<11> out<12> net24 rst rst' vdd vss tff_st_ar
    Xi12 out<7> out<8> net31 rst rst' vdd vss tff_st_ar
    Xi11 out<8> out<9> net38 rst rst' vdd vss tff_st_ar
    Xi10 out<9> out<10> net45 rst rst' vdd vss tff_st_ar
    Xi9 out<10> out<11> net52 rst rst' vdd vss tff_st_ar
    Xi8 out<6> out<7> net59 rst rst' vdd vss tff_st_ar
    Xi7 out<5> out<6> net66 rst rst' vdd vss tff_st_ar
    Xi6 out<4> out<5> net73 rst rst' vdd vss tff_st_ar
    Xi4 out<2> out<3> net87 rst rst' vdd vss tff_st_ar
    Xi3 out<1> out<2> net94 rst rst' vdd vss tff_st_ar
    Xi2 out<0> out<1> net101 rst rst' vdd vss tff_st_ar
    Xi1 rand_in out<0> net108 rst rst' vdd vss tff_st_ar
    Xi5 out<3> out<4> net80 rst rst' vdd vss tff_st_ar
.ENDS
